
** Library name: schem
** Cell name: nand3
** View name: schematic
.subckt nand3 a b c y
m10 net9 c 0 0 nmos L=nl W=nw M=nm
m9 net5 b net9 0 nmos L=nl W=nw M=nm
m1 y a net5 0 nmos L=nl W=nw M=nm
m7 y c vdd! vdd! pmos L=pl W=pw M=pm
m6 y b vdd! vdd! pmos L=pl W=pw M=pm
m0 y a vdd! vdd! pmos L=pl W=pw M=pm
.ends nand3
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_01 a y
m1 y a vdd! vdd! pmos L=2 W=71 M=1
m2 y a 0 0 nmos L=2 W=12 M=1
.ends inv_pcell_01
** End of subcircuit definition.

** Library name: schem
** Cell name: predecode_24
** View name: schematic
.subckt predecode_24 address0 address255 ck inv1 inv1_255
xi36 ck vdd! address0 nand1 nand3 nl=2 nw=9 nm=1 pl=2 pw=3 pm=1
xi37 ck 0 address0 net22 nand3 nl=2 nw=9 nm=1 pl=2 pw=3 pm=1
xi38 ck vdd! address255 nand1_1 nand3 nl=2 nw=9 nm=1 pl=2 pw=3 pm=1
xi39 ck 0 address255 net14 nand3 nl=2 nw=9 nm=1 pl=2 pw=3 pm=1
xu3 net14 net6 inv_pcell_01
xu2 nand1_1 inv1_255 inv_pcell_01
xu1 net22 net10 inv_pcell_01
xu0 nand1 inv1 inv_pcell_01
.ends predecode_24
** End of subcircuit definition.

** Library name: ee313
** Cell name: nor
** View name: schematic
.subckt nor_pcell_2 a b y
m1 mid_a b vdd! vdd! pmos L=2 W=1143 M=1
m2 y a mid_a vdd! pmos L=2 W=1143 M=1
m3 y a 0 0 nmos L=2 W=29 M=1
m4 y b 0 0 nmos L=2 W=400 M=1
.ends nor_pcell_2
** End of subcircuit definition.

** Library name: ee313
** Cell name: nand
** View name: schematic
.subckt nand_pcell_3 a b y
m2 y b vdd! vdd! pmos L=2 W=42 M=15
m0 y a vdd! vdd! pmos L=2 W=42 M=15
m3 mid_a b 0 0 nmos L=2 W=119 M=15
m1 y a mid_a 0 nmos L=2 W=119 M=15
.ends nand_pcell_3
** End of subcircuit definition.

** Library name: ee313
** Cell name: nand
** View name: schematic
.subckt nand_pcell_4 a b y
m2 y b vdd! vdd! pmos L=2 W=42 M=1
m0 y a vdd! vdd! pmos L=2 W=42 M=1
m3 mid_a b 0 0 nmos L=2 W=119 M=1
m1 y a mid_a 0 nmos L=2 W=119 M=1
.ends nand_pcell_4
** End of subcircuit definition.

** Library name: ee313
** Cell name: nor
** View name: schematic
.subckt nor_pcell_5 a b y
m1 mid_a b vdd! vdd! pmos L=2 W=1143 M=15
m2 y a mid_a vdd! pmos L=2 W=1143 M=15
m3 y a 0 0 nmos L=2 W=29 M=15
m4 y b 0 0 nmos L=2 W=400 M=15
.ends nor_pcell_5
** End of subcircuit definition.

** Library name: schem
** Cell name: decode_stage
** View name: schematic
.subckt decode_stage wl0 wl255 predec predec_255 sae sae_b0 sae_b255
xu7 net11 wl_pulldown255 wl255 nor_pcell_2
xu5 net17 wl_pulldown0 wl0 nor_pcell_2
xu1 0 predec net14 nand_pcell_3
xu3 0 predec_255 net8 nand_pcell_3
xu2 vdd! predec_255 net11 nand_pcell_4
xu0 vdd! predec net17 nand_pcell_4
xu6 net14 0 net26 nor_pcell_5
xu8 net8 0 net22 nor_pcell_5
xu9 sae wl0 wl_pulldown0 sae_b0 sae_inv_chain
xu10 sae wl255 wl_pulldown255 sae_b255 sae_inv_chain
.ends decode_stage
** End of subcircuit definition.

** Library name: ee313
** Cell name: nand
** View name: schematic
.subckt nand_pcell_6 a b c y
m2 y b vdd! vdd! pmos L=2 W=20 M=1
m0 y a vdd! vdd! pmos L=2 W=20 M=1
m6 y c vdd! vdd! pmos L=2 W=20 M=1
m3 mid_a b 0 0 nmos L=2 W=74 M=1
m4 mid_b a mid_a 0 nmos L=2 W=74 M=1
m5 y c mid_b 0 nmos L=2 W=74 M=1
.ends nand_pcell_6
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_78 a y
m1 y a vdd! vdd! pmos L=2 W=555 M=1
m2 y a 0 0 nmos L=2 W=92 M=1
.ends inv_pcell_78
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_910 a y
m1 y a vdd! vdd! pmos L=2 W=42 M=1
m2 y a 0 0 nmos L=2 W=119 M=1
.ends inv_pcell_910
** End of subcircuit definition.

** Library name: ee313
** Cell name: nand
** View name: schematic
.subckt nand_pcell_11 a b c y
m2 y b vdd! vdd! pmos L=2 W=20 M=3
m0 y a vdd! vdd! pmos L=2 W=20 M=3
m4 y c vdd! vdd! pmos L=2 W=20 M=3
m3 mid_a b 0 0 nmos L=2 W=74 M=3
m1 mid_b a mid_a 0 nmos L=2 W=74 M=3
m5 y c mid_b 0 nmos L=2 W=74 M=3
.ends nand_pcell_11
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_1213 a y
m1 y a vdd! vdd! pmos L=2 W=42 M=3
m2 y a 0 0 nmos L=2 W=119 M=3
.ends inv_pcell_1213
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_1415 a y
m1 y a vdd! vdd! pmos L=2 W=555 M=3
m2 y a 0 0 nmos L=2 W=92 M=3
.ends inv_pcell_1415
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_16 a y
m1 y a vdd! vdd! pmos L=2 W=1143 M=1
m2 y a 0 0 nmos L=2 W=29 M=1
.ends inv_pcell_16
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_17 a y
m1 y a vdd! vdd! pmos L=2 W=1143 M=3
m2 y a 0 0 nmos L=2 W=29 M=3
.ends inv_pcell_17
** End of subcircuit definition.

** Library name: schem
** Cell name: predecode_416
** View name: schematic
.subckt predecode_416 inv1 inv1_255 predec predec_255 sae_b0 sae_b255
xi17 vdd! inv1_255 sae_b255 net057 nand_pcell_6
xi15 vdd! inv1 sae_b0 net77 nand_pcell_6
xu2 net057 predec_255 inv_pcell_78
xu0 net77 predec inv_pcell_78
xi16 0 inv1 sae_b0 net55 nand_pcell_11
xi18 0 inv1_255 sae_b255 net63 nand_pcell_11
xu1 net55 net69 inv_pcell_1415
xu3 net63 net73 inv_pcell_1415
.ends predecode_416
** End of subcircuit definition.


.subckt sae_inv_chain sae wl wl_pulldown sae_b
x123 sae wl net_sae_1 nand2_1240
x124 net_sae_1 net_sae_2 inv_1241
x125 net_sae_2 sae_b inv_1242
x126 sae_b wl_pulldown inv_1243
.ends sae_inv_chain

.subckt nand2_1240 a b y
m2 y b vdd! vdd! pmos L=2 W=1 M=1
m0 y a vdd! vdd! pmos L=2 W=1 M=1
m3 mid_a b 0 0 nmos L=2 W=3 M=1
m1 y a mid_a 0 nmos L=2 W=3 M=1
.ends nand2_1240

.subckt inv_1241 a y
m1 y a vdd! vdd! pmos L=2 W=19 M=1
m2 y a 0 0 nmos L=2 W=3 M=1
.ends inv_1241

.subckt inv_1242 a y
m1 y a vdd! vdd! pmos L=2 W=23 M=1
m2 y a 0 0 nmos L=2 W=47 M=1
.ends inv_1242

.subckt inv_1243 a y
m1 y a vdd! vdd! pmos L=2 W=436 M=1
m2 y a 0 0 nmos L=2 W=73 M=1
.ends inv_1243
