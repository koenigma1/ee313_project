
** Library name: project_2012_part1_sol
** Cell name: task3
** View name: schematic
xcbl bl0 bl_b0 wl255 vdd gnd 0 vdd! mc m=1
xi5 net57 net56 wl255 vdd gnd 0 vdd! mc m=254
xcbr bl63 bl_b63 wl255 vdd gnd 0 vdd! mc m=1
xi4 bl63 bl_b63 0 vdd gnd 0 vdd! mc m=254
xi3 net57 net56 0 vdd gnd 0 vdd! mc m=64.516e3
xi2 bl0 bl_b0 0 vdd gnd 0 vdd! mc m=254
xctr bl63 bl_b63 wl0 vdd gnd 0 vdd! mc m=1
xi1 net57 net56 wl0 vdd gnd 0 vdd! mc m=254
xctl bl0 bl_b0 wl0 vdd gnd 0 vdd! mc m=1
xwritel bl0 bl_b0 blpc_b vdd! 0 0 vdd! write m=1
xwritem net57 net56 blpc_b vdd! 0 0 vdd! write m=254
xwriter bl63 bl_b63 blpc_b vdd! 0 0 vdd! write m=1
xi17 wl0 wl255 a0 a255 ck decoder_schematic
