
** Library name: schem
** Cell name: nand3
** View name: schematic
.subckt nand3 a b c y
m10 net9 c 0 0 nmos L=nl W=nw M=nm
m9 net5 b net9 0 nmos L=nl W=nw M=nm
m1 y a net5 0 nmos L=nl W=nw M=nm
m7 y c vdd! vdd! pmos L=pl W=pw M=pm
m6 y b vdd! vdd! pmos L=pl W=pw M=pm
m0 y a vdd! vdd! pmos L=pl W=pw M=pm
.ends nand3
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_0 a y
m1 y a vdd! vdd! pmos L=2 W=41 M=1
m2 y a 0 0 nmos L=2 W=7 M=1
.ends inv_pcell_0
** End of subcircuit definition.

** Library name: schem
** Cell name: predecode_24
** View name: schematic
.subckt predecode_24 address0 address255 ck inv1 inv1_255
xi36 ck vdd! address0 nand1 nand3 nl=2 nw=9 nm=1 pl=2 pw=3 pm=1
xi37 ck 0 address0 net22 nand3 nl=2 nw=9 nm=1 pl=2 pw=3 pm=1
xi38 ck vdd! address255 nand1_1 nand3 nl=2 nw=9 nm=1 pl=2 pw=3 pm=1
xi39 ck 0 address255 net14 nand3 nl=2 nw=9 nm=1 pl=2 pw=3 pm=1
xu3 net14 net6 inv_pcell_0
xu2 nand1_1 inv1_255 inv_pcell_0
xu1 net22 net10 inv_pcell_0
xu0 nand1 inv1 inv_pcell_0
.ends predecode_24
** End of subcircuit definition.

** Library name: ee313
** Cell name: nand
** View name: schematic
.subckt nand_pcell_1 a b y
m2 y b vdd! vdd! pmos L=2 W=340 M=1
m0 y a vdd! vdd! pmos L=2 W=340 M=1
m3 mid_a b 0 0 nmos L=2 W=57 M=1
m1 y a mid_a 0 nmos L=2 W=57 M=1
.ends nand_pcell_1
** End of subcircuit definition.

** Library name: ee313
** Cell name: nand
** View name: schematic
.subckt nand_pcell_2 a b y
m2 y b vdd! vdd! pmos L=2 W=340 M=15
m0 y a vdd! vdd! pmos L=2 W=340 M=15
m3 mid_a b 0 0 nmos L=2 W=57 M=15
m1 y a mid_a 0 nmos L=2 W=57 M=15
.ends nand_pcell_2
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_3 a y
m1 y a vdd! vdd! pmos L=2 W=292 M=1
m2 y a 0 0 nmos L=2 W=583 M=1
.ends inv_pcell_3
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_4 a y
m1 y a vdd! vdd! pmos L=2 W=292 M=15
m2 y a 0 0 nmos L=2 W=583 M=15
.ends inv_pcell_4
** End of subcircuit definition.

** Library name: schem
** Cell name: decode_stage
** View name: schematic
.subckt decode_stage wl0 wl255 predec predec_255
xu2 vdd! predec_255 net11 nand_pcell_1
xu0 vdd! predec net17 nand_pcell_1
xu3 0 predec_255 net8 nand_pcell_2
xu1 0 predec net14 nand_pcell_2
xu7 net11 wl255 inv_pcell_3
xu5 net17 wl0 inv_pcell_3
xu8 net8 net22 inv_pcell_4
xu6 net14 net26 inv_pcell_4
.ends decode_stage
** End of subcircuit definition.

** Library name: ee313
** Cell name: nand
** View name: schematic
.subckt nand_pcell_5 a b y
m2 y b vdd! vdd! pmos L=2 W=34 M=1
m0 y a vdd! vdd! pmos L=2 W=34 M=1
m3 mid_a b 0 0 nmos L=2 W=6 M=1
m1 y a mid_a 0 nmos L=2 W=6 M=1
.ends nand_pcell_5
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_6 a y
m1 y a vdd! vdd! pmos L=2 W=31 M=1
m2 y a 0 0 nmos L=2 W=62 M=1
.ends inv_pcell_6
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_7 a y
m1 y a vdd! vdd! pmos L=2 W=31 M=3
m2 y a 0 0 nmos L=2 W=62 M=3
.ends inv_pcell_7
** End of subcircuit definition.

** Library name: ee313
** Cell name: nand
** View name: schematic
.subckt nand_pcell_8 a b y
m2 y b vdd! vdd! pmos L=2 W=34 M=3
m0 y a vdd! vdd! pmos L=2 W=34 M=3
m3 mid_a b 0 0 nmos L=2 W=6 M=3
m1 y a mid_a 0 nmos L=2 W=6 M=3
.ends nand_pcell_8
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_9 a y
m1 y a vdd! vdd! pmos L=2 W=444 M=1
m2 y a 0 0 nmos L=2 W=74 M=1
.ends inv_pcell_9
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_10 a y
m1 y a vdd! vdd! pmos L=2 W=410 M=1
m2 y a 0 0 nmos L=2 W=820 M=1
.ends inv_pcell_10
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_11 a y
m1 y a vdd! vdd! pmos L=2 W=444 M=3
m2 y a 0 0 nmos L=2 W=74 M=3
.ends inv_pcell_11
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_12 a y
m1 y a vdd! vdd! pmos L=2 W=410 M=3
m2 y a 0 0 nmos L=2 W=820 M=3
.ends inv_pcell_12
** End of subcircuit definition.

** Library name: schem
** Cell name: predecode_416
** View name: schematic
.subckt predecode_416 inv1 inv1_255 predec predec_255
xi15 vdd! inv1 net77 nand_pcell_5
xi17 vdd! inv1_255 net057 nand_pcell_5
xu0 net77 net032 inv_pcell_6
xu2 net057 net036 inv_pcell_6
xu1 net55 net69 inv_pcell_7
xu3 net63 net73 inv_pcell_7
xi16 0 inv1 net55 nand_pcell_8
xi18 0 inv1_255 net63 nand_pcell_8
xu15 net032 net046 inv_pcell_9
xu13 net036 net052 inv_pcell_9
xu10 net052 predec_255 inv_pcell_10
xu8 net046 predec inv_pcell_10
xu14 net69 net049 inv_pcell_11
xu12 net73 net043 inv_pcell_11
xu11 net043 net024 inv_pcell_12
xu9 net049 net028 inv_pcell_12
.ends predecode_416
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_13 a y
m1 y a vdd! vdd! pmos L=2 W=8
m2 y a 0 0 nmos L=2 W=4
.ends inv_pcell_13
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_14 a y
m1 y a vdd! vdd! pmos L=2 W=12
m2 y a 0 0 nmos L=2 W=24
.ends inv_pcell_14
** End of subcircuit definition.

** Library name: schem
** Cell name: write
** View name: schematic
.subckt write bl0 bl_b0 blpc_b wrdata wren0 inh_bulk_n inh_bulk_p
m5 bl0 blpc_b vdd! inh_bulk_p pmos L=2 W=80
m1 bl0 blpc_b bl_b0 inh_bulk_p pmos L=2 W=80
m0 bl_b0 blpc_b vdd! inh_bulk_p pmos L=2 W=80
m4 net23 wren0 bl_b0 inh_bulk_n nmos L=2 W=90
m3 net26 wren0 bl0 inh_bulk_n nmos L=2 W=90
xu0 wrdata net18 inv_pcell_13
xu2 wrdata net23 inv_pcell_14
xu1 net18 net26 inv_pcell_14
.ends write
** End of subcircuit definition.

** Library name: schem
** Cell name: mc
** View name: schematic
.subckt mc bl bl_b wl vdd vss inh_bulk_n inh_bulk_p
m5 bit bit_b vss inh_bulk_n nmos L=2 W=6
m4 bit_b bit vss inh_bulk_n nmos L=2 W=6
m1 bl_b wl bit_b inh_bulk_n nmos L=2 W=4
m0 bl wl bit inh_bulk_n nmos L=2 W=4
m2 bit_b bit vdd inh_bulk_p pmos L=2 W=4
m3 bit bit_b vdd inh_bulk_p pmos L=2 W=4
c2 bl 0 88e-18
c1 bl_b 0 88e-18
c0 wl 0 140e-18
.ends mc
** End of subcircuit definition.

** Library name: schem
** Cell name: SRAM
** View name: schematic
.subckt SRAM bl0 bl63 bl_b0 bl_b63 blpc_b wl0 wl255 inh_bulk_n inh_bulk_p
xi16 bl63 bl_b63 blpc_b vdd! 0 inh_bulk_n inh_bulk_p write m=1
xi17 net9 net8 blpc_b vdd! 0 inh_bulk_n inh_bulk_p write m=254
xi14 bl0 bl_b0 blpc_b vdd! 0 inh_bulk_n inh_bulk_p write m=1
xiBOTTOM_RIGHT bl63 bl_b63 wl255 vdd! gnd inh_bulk_n inh_bulk_p mc m=1
xi13 net9 net8 wl255 vdd! gnd inh_bulk_n inh_bulk_p mc m=254
xiBOTTOM_LEFT bl0 bl_b0 wl255 vdd! gnd inh_bulk_n inh_bulk_p mc m=1
xi11 bl0 bl_b0 0 vdd! gnd inh_bulk_n inh_bulk_p mc m=254
xi10 net9 net8 0 vdd! gnd inh_bulk_n inh_bulk_p mc m=64.52e3
xi12 bl63 bl_b63 0 vdd! gnd inh_bulk_n inh_bulk_p mc m=254
xiTOP_RIGHT bl63 bl_b63 wl0 vdd! gnd inh_bulk_n inh_bulk_p mc m=1
xi9 net9 net8 wl0 vdd! gnd inh_bulk_n inh_bulk_p mc m=254
xiTOP_LEFT bl0 bl_b0 wl0 vdd! gnd inh_bulk_n inh_bulk_p mc m=1
.ends SRAM
** End of subcircuit definition.

** Library name: schem
** Cell name: task3
** View name: schematic
xi5 address0 address255 ck net2 net1 predecode_24
xi4 net2 net1 net14 net17 predecode_416
xi1 wl0 wl255 net14 net17 decode_stage
c_sideload2 net17 0 22.53e-15
c_sideload net14 0 22.53e-15
xiSRAM bl0 bl63 bl_b0 bl_b63 blpc_b wl0 wl255 0 vdd! SRAM
