
** Library name: Proyect
** Cell name: mc
** View name: schematic
.subckt mc bl bl_b wl vdd vss inh_bulk_n inh_bulk_p
m5 bit bit_b vss inh_bulk_n nmos L=2 W=6
m4 bit_b bit vss inh_bulk_n nmos L=2 W=6
m1 bl_b wl bit_b inh_bulk_n nmos L=2 W=4
m0 bl wl bit inh_bulk_n nmos L=2 W=4
m2 bit_b bit vdd inh_bulk_p pmos L=2 W=4
m3 bit bit_b vdd inh_bulk_p pmos L=2 W=4
c2 bl 0 88e-18
c1 bl_b 0 88e-18
c0 wl 0 140e-18
.ends mc
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_0 a y
m1 y a vdd! vdd! pmos L=2 W=8
m2 y a 0 0 nmos L=2 W=4
.ends inv_pcell_0
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_1 a y
m1 y a vdd! vdd! pmos L=2 W=12
m2 y a 0 0 nmos L=2 W=24
.ends inv_pcell_1
** End of subcircuit definition.

** Library name: Proyect
** Cell name: write
** View name: schematic
.subckt write bl0 bl_b0 blpc_b wrdata wren0 inh_bulk_n inh_bulk_p
m5 bl0 blpc_b vdd! inh_bulk_p pmos L=2 W=80
m1 bl0 blpc_b bl_b0 inh_bulk_p pmos L=2 W=80
m0 bl_b0 blpc_b vdd! inh_bulk_p pmos L=2 W=80
m4 net23 wren0 bl_b0 inh_bulk_n nmos L=2 W=90
m3 net26 wren0 bl0 inh_bulk_n nmos L=2 W=90
xu0 wrdata net18 inv_pcell_0
xu2 wrdata net23 inv_pcell_1
xu1 net18 net26 inv_pcell_1
.ends write
** End of subcircuit definition.

** Library name: Proyect
** Cell name: SRAM
** View name: schematic
xi8 bl63 bl_b63 wl255 vdd! gnd 0 vdd! mc m=1
xi13 net9 net8 wl255 vdd! gnd 0 vdd! mc m=254
xi6 bl0 bl_b0 wl255 vdd! gnd 0 vdd! mc m=1
xi11 bl0 bl_b0 0 vdd! gnd 0 vdd! mc m=254
xi10 net9 net8 0 vdd! gnd 0 vdd! mc m=64.516e3
xi12 bl63 bl_b63 0 vdd! gnd 0 vdd! mc m=254
xi2 bl63 bl_b63 wl0 vdd! gnd 0 vdd! mc m=1
xi9 net9 net8 wl0 vdd! gnd 0 vdd! mc m=254
xi0 bl0 bl_b0 wl0 vdd! gnd 0 vdd! mc m=1
xi16 bl63 bl_b63 blpc_b vdd! 0 0 vdd! write m=1
xi17 net9 net8 blpc_b vdd! 0 0 vdd! write m=254
xi14 bl0 bl_b0 blpc_b vdd! 0 0 vdd! write m=1
