
** Library name: Proyect
** Cell name: mc
** View name: schematic
.subckt mc bl bl_b wl vdd vss inh_bulk_n inh_bulk_p
m5 bit bit_b vss inh_bulk_n nmos L=2 W=6
m4 bit_b bit vss inh_bulk_n nmos L=2 W=6
m1 bl_b wl bit_b inh_bulk_n nmos L=2 W=4
m0 bl wl bit inh_bulk_n nmos L=2 W=4
m2 bit_b bit vdd inh_bulk_p pmos L=2 W=4
m3 bit bit_b vdd inh_bulk_p pmos L=2 W=4
c2 bl 0 88e-18
c1 bl_b 0 88e-18
c0 wl 0 140e-18
.ends mc
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_0 a y
m1 y a vdd! vdd! pmos L=2 W=8
m2 y a 0 0 nmos L=2 W=4
.ends inv_pcell_0
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt inv_pcell_1 a y
m1 y a vdd! vdd! pmos L=2 W=12
m2 y a 0 0 nmos L=2 W=24
.ends inv_pcell_1
** End of subcircuit definition.

** Library name: Proyect
** Cell name: write
** View name: schematic
.subckt write bl0 bl_b0 blpc_b wrdata wren0 inh_bulk_n inh_bulk_p
Vbl bl0 bl0_prime dc 0
m2 bl0_prime blpc_b vdd! inh_bulk_p pmos L=2 W=80
m1 bl0_prime blpc_b bl_b0 inh_bulk_p pmos L=2 W=80
m0 bl_b0 blpc_b vdd! inh_bulk_p pmos L=2 W=80
m4 net23 wren0 bl_b0 inh_bulk_n nmos L=2 W=90
m3 net26 wren0 bl0_prime inh_bulk_n nmos L=2 W=90
xu0 wrdata net18 inv_pcell_0
xu2 wrdata net23 inv_pcell_1
xu1 net18 net26 inv_pcell_1
.ends write
** End of subcircuit definition.

******************************
** SENSE AMP POSTED HERE

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt sense_inv_pcell_0 a y
m1 y a vdd! vdd! pmos L=2 W=24
m2 y a 0 0 nmos L=2 W=12
.ends sense_inv_pcell_0
** End of subcircuit definition.

** Library name: ee313
** Cell name: inv
** View name: schematic
.subckt sense_inv_pcell_1 a y
m1 y a vdd! vdd! pmos L=2 W=100
m2 y a 0 0 nmos L=2 W=50
.ends sense_inv_pcell_1
** End of subcircuit definition.

** Library name: schem
** Cell name: sense
** View name: schematic
.subckt sense bl0 bl_b0 sel_b0 sapc_b sae out out_b  
m4 sbl_b sbl vdd! vdd! pmos L=2 W=4
m3 vdd! sbl_b sbl vdd! pmos L=2 W=4
meq sbl sapc_b sbl_b vdd! pmos L=2 W=8
mpc2 vdd! sapc_b sbl_b vdd! pmos L=2 W=8
mpc sbl sapc_b vdd! vdd! pmos L=2 W=8
miso_b sbl_b sae cmbl_b vdd! pmos L=2 W=12
miso sbl sae cmbl vdd! pmos L=2 W=12
mmx4_b cmbl_b vdd! vdd! vdd! pmos L=2 W=24
mmx4 cmbl vdd! vdd! vdd! pmos L=2 W=24
mmx3_b cmbl_b vdd! vdd! vdd! pmos L=2 W=24
mmx3 cmbl vdd! vdd! vdd! pmos L=2 W=24
mmx2_b cmbl_b vdd! vdd! vdd! pmos L=2 W=24
mmx2 cmbl vdd! vdd! vdd! pmos L=2 W=24
mmx_b cmbl_b sel_b0 bl_b0 vdd! pmos L=2 W=24
mmx cmbl sel_b0 bl0 vdd! pmos L=2 W=24
mtail tail sae 0 0 nmos L=2 W=8
m1 tail sbl_b sbl 0 nmos L=2 W=6
m2 sbl_b sbl tail 0 nmos L=2 W=6
c1 sapc_b 0 560e-18
c0 sae 0 560e-18
xu1 sbl_b out sense_inv_pcell_0
xu0 sbl out_b sense_inv_pcell_0
xu3 out net70 sense_inv_pcell_1
xu2 out_b net71 sense_inv_pcell_1
.ends
******************************

** Library name: Proyect
** Cell name: SRAM
** View name: schematic
xi8 bl63 bl_b63 wl255 vdd! gnd 0 vdd! mc m=1
xi13 net9 net8 wl255 vdd! gnd 0 vdd! mc m=254
xi6 bl0 bl_b0 wl255 vdd! gnd 0 vdd! mc m=1
xi11 bl0 bl_b0 0 vdd! gnd 0 vdd! mc m=254
xi10 net9 net8 0 vdd! gnd 0 vdd! mc m=64.516e3
xi12 bl63 bl_b63 0 vdd! gnd 0 vdd! mc m=254
xi2 bl63 bl_b63 wl0 vdd! gnd 0 vdd! mc m=1
xi9 net9 net8 wl0 vdd! gnd 0 vdd! mc m=254
xiTOP_LEFT bl0 bl_b0 wl0 vdd! gnd 0 vdd! mc m=1
xi16 bl63 bl_b63 blpc_b vdd! 0 0 vdd! write m=1
xi17 net9 net8 blpc_b vdd! 0 0 vdd! write m=254
xi14 bl0 bl_b0 blpc_b vdd! 0 0 vdd! write m=1
xsense bl_0 bl_b0 0 sapc_b sae out out_b sense

